module tb();
logic [3:0]d[7:0];
logic [3:0]y;
logic [2:0]s;

d[0]=3'b1000;
d[1]=3'b1001;
d[2]=3'b1010;
d[3]=3'b1011;
d[4]=3'b1100;
d[5]=3'b1101;
d[6]=3'b1110;
d[7]=3'b1111;

mux81 m1(d,s,y);
initial begin
s[0]=0;s[1]=0;s[2]=0;
#10
s[0]=0;s[1]=0;s[2]=1;
#10
s[0]=0;s[1]=1;s[2]=0;
#10
s[0]=0;s[1]=1;s[2]=1;
#10
s[0]=1;s[1]=0;s[2]=0;
#10
s[0]=1;s[1]=0;s[2]=1;
#10
s[0]=1;s[1]=1;s[2]=0;
#10
s[0]=1;s[1]=1;s[2]=1;
end 
endmodule
